LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY fpAdd_Controller IS
  port( Mantissa_Overflow : IN std_logic; 
    LargerB : OUT std_logic);
END fpAdd_Controller;

ARCHITECTURE struct OF fpAdd_Controller IS
BEGIN
  
END struct;